library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MIPS is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC);
end MIPS;

architecture Behavioral of MIPS is

begin


end Behavioral;

